/home/01fe21bee114/internship/DFT_LIB/LEF/FreePDK45_lib_v1.0.MOD.lef