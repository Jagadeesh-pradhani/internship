/home/01fe21bee114/internship/DFT_LIB/LEF/NanGate_15nm_OCL.tech.lef