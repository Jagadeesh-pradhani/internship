/home/01fe21bee114/internship/DFT_LIB/LIB/slow.vhd